`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:03:08 04/13/2012 
// Design Name: 
// Module Name:    dispatcher 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dispatcher(
    input [4:0] a1,
    input [4:0] a2,
    input [4:0] a3,
    input [4:0] a4
    );


endmodule
