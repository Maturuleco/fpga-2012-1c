`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    11:09:47 04/13/2012 
// Design Name: 
// Module Name:    dilplay_cont 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module dilplay_cont(
	 input wire clk,
    input wire tick,
	 input wire reset,
    input wire en,
    input wire up,
    input wire[3:0] d,
    input wire syn_clr,
    input wire load,
    output wire max_tick,
    output wire min_tick,
    output wire [7:0] sseg,
	 output [3:0] an
    );
	 
	wire[3:0] q;
	wire tick_damped;
	db_fsm antiruido (
		.clk(clk),
		.reset(reset),
		.sw(tick),
		.db(tick_damped)
	);
	universal_bin_count_4bit  ubc (
		.clk(tick_damped),
		.reset(reset),
		.en(en),
		.up(up),
		.d(d),
		.syn_clr(syn_clr),
		.load(load),
		.max_tick(max_tick),
		.min_tick(min_tick),
		.q(q)
	);
	
	wire [3:0] s1, s2, s3;
	wire [7:0] salida1, salida2, salida3;

	bit_to_3hexa_digits	refactor	( .entrada(q), .h1(s1), .h2(s2), .h3(s3) );

	hex_to_sseg	numero1	(.hex(s1), .dp(1'b0), .sseg(salida1));
	hex_to_sseg	numero2	(.hex(s2), .dp(1'b0), .sseg(salida2));
	hex_to_sseg	numero3	(.hex(s3), .dp(1'b0), .sseg(salida3));
	
	disp_mux		display	(.in0(salida1), .in1(salida2), .in2(salida3), .in3(1), .an(an), .sseg(sseg), .clk(clk), .reset(reset) );

endmodule
